library verilog;
use verilog.vl_types.all;
entity sumador_completo_vlg_check_tst is
    port(
        o_count         : in     vl_logic;
        o_f             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end sumador_completo_vlg_check_tst;
