library verilog;
use verilog.vl_types.all;
entity ejercicio1_diagram_block_vlg_vec_tst is
end ejercicio1_diagram_block_vlg_vec_tst;
