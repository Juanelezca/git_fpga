library verilog;
use verilog.vl_types.all;
entity ejercicio1_vlg_vec_tst is
end ejercicio1_vlg_vec_tst;
