library verilog;
use verilog.vl_types.all;
entity ejercicio1_diagram_block_vlg_check_tst is
    port(
        LED             : in     vl_logic;
        LED8            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end ejercicio1_diagram_block_vlg_check_tst;
